/***********************************************module and port declartion*************************************************/
module reset_synchronizer_deasertion (
input wire clk,rst,
output reg reset_senchronizer
);
/**************************************************************************************************************************/

/***********************************************signal declartion**********************************************************/        
reg sign;
reg D;
assign D = 1;
/**************************************************************************************************************************/

/**************************************************************************************************************************/
always@(posedge clk or negedge rst)
begin
sign <= D  ;
reset_senchronizer <= sign ;
end
endmodule
/**************************************************************************************************************************/